-- Vhdl test bench created from schematic C:\Users\Seres\Desktop\DIGIT\digit_remake\knight_rider_remake\kr_remake.sch - Fri Nov 22 15:01:05 2019
--
-- Notes: 
-- 1) This testbench template has been automatically generated using types
-- std_logic and std_logic_vector for the ports of the unit under test.
-- Xilinx recommends that these types always be used for the top-level
-- I/O of a design in order to guarantee that the testbench will bind
-- correctly to the timing (post-route) simulation model.
-- 2) To use this template as your testbench, change the filename to any
-- name of your choice with the extension .vhd, and use the "Source->Add"
-- menu in Project Navigator to import the testbench. Then
-- edit the user defined section below, adding code to generate the 
-- stimulus for your design.
--
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;
LIBRARY UNISIM;
USE UNISIM.Vcomponents.ALL;
ENTITY kr_remake_kr_remake_sch_tb IS
END kr_remake_kr_remake_sch_tb;
ARCHITECTURE behavioral OF kr_remake_kr_remake_sch_tb IS 

   COMPONENT kr_remake
   PORT( q	:	OUT	STD_LOGIC_VECTOR (3 DOWNTO 0); 
          en	:	IN	STD_LOGIC; 
          clk	:	IN	STD_LOGIC);
   END COMPONENT;

   SIGNAL q	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
   SIGNAL en	:	STD_LOGIC;
   SIGNAL clk	:	STD_LOGIC;

BEGIN

   UUT: kr_remake PORT MAP(
		q => q, 
		en => en, 
		clk => clk
   );

-- *** Test Bench - User Defined Section ***
   tb : PROCESS
   BEGIN
	   en <= '1';
		clk <= '0';
		wait for 4 us;
		clk <= '1';
		wait for 4 us;
   END PROCESS;
-- *** End Test Bench - User Defined Section ***

END;
