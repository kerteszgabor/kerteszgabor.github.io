-- Vhdl test bench created from schematic C:\Users\Seres\Desktop\DIGIT\digit_remake\szamlalo3_remake\szamlalo3_remake.sch - Fri Nov 22 15:28:10 2019
--
-- Notes: 
-- 1) This testbench template has been automatically generated using types
-- std_logic and std_logic_vector for the ports of the unit under test.
-- Xilinx recommends that these types always be used for the top-level
-- I/O of a design in order to guarantee that the testbench will bind
-- correctly to the timing (post-route) simulation model.
-- 2) To use this template as your testbench, change the filename to any
-- name of your choice with the extension .vhd, and use the "Source->Add"
-- menu in Project Navigator to import the testbench. Then
-- edit the user defined section below, adding code to generate the 
-- stimulus for your design.
--
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;
LIBRARY UNISIM;
USE UNISIM.Vcomponents.ALL;
ENTITY szamlalo3_remake_szamlalo3_remake_sch_tb IS
END szamlalo3_remake_szamlalo3_remake_sch_tb;
ARCHITECTURE behavioral OF szamlalo3_remake_szamlalo3_remake_sch_tb IS 

   COMPONENT szamlalo3_remake
   PORT( sw	:	IN	STD_LOGIC; 
          clk	:	IN	STD_LOGIC; 
          q	:	OUT	STD_LOGIC_VECTOR (3 DOWNTO 0));
   END COMPONENT;

   SIGNAL sw	:	STD_LOGIC;
   SIGNAL clk	:	STD_LOGIC;
   SIGNAL q	:	STD_LOGIC_VECTOR (3 DOWNTO 0);

BEGIN

   UUT: szamlalo3_remake PORT MAP(
		sw => sw, 
		clk => clk, 
		q => q
   );

-- *** Test Bench - User Defined Section ***
   tb : PROCESS
   BEGIN
     sw <= '1';
	  clk <= '0';
	  wait for 4 us;
	  clk <= '1';
	  wait for 4 us;
   END PROCESS;
-- *** End Test Bench - User Defined Section ***

END;
